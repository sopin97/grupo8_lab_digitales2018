// RAM_WIDTH -> tama;o de una palabra
// RAM_HEIGHT -> numero de "slots" en la RAM
module RAM_reader #(parameter RAM_WIDTH = 8, parameter RAM_DEPTH = (1024*768*3*8)/RAM_WIDTH)
(
  input logic [RAM_WIDTH-1:0] data,
  input logic rst, clk, refresh_data,
  output logic [ADRESS_BITS-1:0] adress,
  output logic [RAM_WIDTH-1:0] data_out
);
  
  localparam ADRESS_BITS = $clog2(RAM_DEPTH); // numero de bits de adress
  logic [ADRESS_BITS-1:0] next_adress;
  
  enum logic [1:0] {IDLE, READ_DATA, REFRESH_ADRESS, WAIT} next_state, state;
  logic [ADRESS_BITS-1:0] next_adress;
  logic [RAM_WIDTH-1:0] next_output;

  always_ff @(posedge clk) begin
    if (rst) begin
      data_out <= 'd0;
      adress <= 'd0;
    else begin
      data_out <= next_output;
      adress <= next_adress;
    end
   end
  always_comb begin
    next_state = state;
    next_output = data_out;
    next_adress = adress;
    case(state)
      IDLE: begin
        if (refresh_data)
          next_state = READ_DATA;
      end
      READ_DATA: begin
        next_output = data;
        next_state = REFRESH_ADRESS;
      end
      REFRESH_ADRESS:
        
        next_adress = adress + 'd1;
        next_state = WAIT;
      WAIT:
        if (!refresh_data)
          next_state = IDLE;
      
  end
  endmodule
