module convertidor (
